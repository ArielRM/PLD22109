
module src_and_probes (
	source,
	probe);	

	output	[3:0]	source;
	input	[2:0]	probe;
endmodule
