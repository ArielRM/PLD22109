
module unnamed (
	probe,
	source);	

	input	[15:0]	probe;
	output	[16:0]	source;
endmodule
